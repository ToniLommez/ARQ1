// -------------------------
// Recuperação 01
// Nome: Marcos Antonio Lommez Candido Ribeiro
// Matricula: 771157
// 31/10/2022
// -------------------------

module A0113 ( output s, input a, input b, input c);
    assign s = ~((~a|~b) & ~(a&c));
endmodule

module questao03;
    reg a, b, c; // Variaveis
    reg contador;
    wire s1;     // Respostas

    A0113 A01131 ( s1, a, b, c );

    initial
        begin: initial_values
            a = 1'b0; b = 1'b0; c = 1'b0; contador = 0;
        end

    initial
        begin: main
            $display ( "\n" );
            $display ( "||==============================================||" );
            $display ( "||        Marcos Antonio Lommez - 771157        ||" );
            $display ( "||==============================================||" );
            $display ( "||       m  0 | 1 | 2 | 3 | 4 | 5 | 6 | 7       ||" );
            $display ( "||          0 | 0 | 0 | 0 | 0 | 1 | 1 | 1       ||" );
            $display ( "||==============================================||" );
            $display ( "||    m    || variaveis || expressao ||  saida  ||" );
            $display ( "||---------||-----------||-----------||---------||" );
            #1 a = 0; b = 0; c = 0; contador = 0;
            #0 $display ( "||    %1d    ||   %b %b %b   || %sa%s.b%s.c%s ||    %b    ||", $time, a, b, c, (s1?">":" "), (a?" ":"'"), (b?" ":"'"), (c?" ":"'"), s1);
            #1 a = 0; b = 0; c = 1; contador = 1;
            #0 $display ( "||    %1d    ||   %b %b %b   || %sa%s.b%s.c%s ||    %b    ||", $time, a, b, c, (s1?">":" "), (a?" ":"'"), (b?" ":"'"), (c?" ":"'"), s1);
            #1 a = 0; b = 1; c = 0; contador = 2;
            #0 $display ( "||    %1d    ||   %b %b %b   || %sa%s.b%s.c%s ||    %b    ||", $time, a, b, c, (s1?">":" "), (a?" ":"'"), (b?" ":"'"), (c?" ":"'"), s1);
            #1 a = 0; b = 1; c = 1; contador = 3;
            #0 $display ( "||    %1d    ||   %b %b %b   || %sa%s.b%s.c%s ||    %b    ||", $time, a, b, c, (s1?">":" "), (a?" ":"'"), (b?" ":"'"), (c?" ":"'"), s1);
            #1 a = 1; b = 0; c = 0; contador = 4;
            #0 $display ( "||    %1d    ||   %b %b %b   || %sa%s.b%s.c%s ||    %b    ||", $time, a, b, c, (s1?">":" "), (a?" ":"'"), (b?" ":"'"), (c?" ":"'"), s1);
            #1 a = 1; b = 0; c = 1; contador = 5;
            #0 $display ( "||    %1d    ||   %b %b %b   || %sa%s.b%s.c%s ||    %b    ||", $time, a, b, c, (s1?">":" "), (a?" ":"'"), (b?" ":"'"), (c?" ":"'"), s1);
            #1 a = 1; b = 1; c = 0; contador = 6;
            #0 $display ( "||    %1d    ||   %b %b %b   || %sa%s.b%s.c%s ||    %b    ||", $time, a, b, c, (s1?">":" "), (a?" ":"'"), (b?" ":"'"), (c?" ":"'"), s1);
            #1 a = 1; b = 1; c = 1; contador = 7;
            #0 $display ( "||    %1d    ||   %b %b %b   || %sa%s.b%s.c%s ||    %b    ||", $time, a, b, c, (s1?">":" "), (a?" ":"'"), (b?" ":"'"), (c?" ":"'"), s1);
            #0 $display ( "||==============================================||" );
            #0 $display ( "||  SoP = (a .b'.c ) + (a .b .c') + (a .b .c )  ||" );
            #0 $display ( "||==============================================||" );
            #1 $display ( "\n" );
        end
endmodule

/* 
||==============================================||
||        Marcos Antonio Lommez - 771157        ||
||==============================================||
||       m  0 | 1 | 2 | 3 | 4 | 5 | 6 | 7       ||
||          0 | 0 | 0 | 0 | 0 | 1 | 1 | 1       ||
||==============================================||
||    m    || variaveis || expressao ||  saida  ||
||---------||-----------||-----------||---------||
||    1    ||   0 0 0   ||  a'.b'.c' ||    0    ||
||    2    ||   0 0 1   ||  a'.b'.c  ||    0    ||
||    3    ||   0 1 0   ||  a'.b .c' ||    0    ||
||    4    ||   0 1 1   ||  a'.b .c  ||    0    ||
||    5    ||   1 0 0   ||  a .b'.c' ||    0    ||
||    6    ||   1 0 1   || >a .b'.c  ||    1    ||
||    7    ||   1 1 0   || >a .b .c' ||    1    ||
||    8    ||   1 1 1   || >a .b .c  ||    1    ||
||==============================================||
||  SoP = (a .b'.c ) + (a .b .c') + (a .b .c )  ||
||==============================================||
 */